// SIN_S11_S11.v
//
//
//M13t          :tiny DBG ifdef switch
//L7Ew          :add CK_EE_i
//KAHs          :add 1dly and mach modern coding rule
//KAFw          :touch port config
//170522su      :debug C_XCLIP_1POINT0
//170516tu      :add EN_CK_i , CK&XARST add tail suffix _i
//               mod  C_1POINT0_ON  -> C_XCLIP_1POINT0
//151220su      :mk easy to inference ROM coding in MAX10
//              :mk easy to inference ROM coding in Cyclone I
//151218fr      : rm ~~~_inc.v
//                sin table +0.5
//                retruct external rom ~~~_inc.v
//151215tu      :mod selectanble to clip 1.0
//151213su      :1st.
`include "../MISC/define.vh"
`ifndef SIN_S11_S11
module SIN_S11_S11
(
      `in`tri1          CK_i  
    , `in`tri1          XARST_i
    , `in`tri1          CK_EE_i 
    , `in`tri0[7:0]     B_IN_DAT_DLYs_i
    , `in`tri0[11:0]    DATs_i     //2's -h800 0 +7FFF
    , `out`w  [11:0]    SINs_o     //2's -h7ff 0 +h7FF
    , `out`w            DONE_o
    , `out`w[7:0]       B_OUT_DAT_DLYs_o
) ;
    localparam C_DAT_DLYs = 1 ;

    // main
    `w down_curve = DATs_i[10] ;
    `w`s[ 9:0] sin_adr_s = ( down_curve ) ? -DATs_i[ 9 :0] : DATs_i[9 :0] ;

    // 3CK_i dly
    `w[ 8:0] SIN_ROM_DATs   ;
    `w[ 7:0] B_ROM_DAT_DLYs ;
    `w       SIN_CODE_DONE  ;
    SIN_ROM_S11_S11
        SIN_ROM_S11_S11
        (     .CK_i             ( CK_i              )
            , .XARST_i          ( XARST_i           )
            , .CK_EE_i          ( CK_EE_i           )
            , .B_IN_DAT_DLYs_i  ( B_IN_DAT_DLYs_i   )
            , .ADRs_i           ( sin_adr_s         )
            , .QQs_o            ( SIN_ROM_DATs      )
            , .DONE_o           ( SIN_CODE_DONE     )
            , .B_OUT_DAT_DLYs_o ( B_ROM_DAT_DLYs    )
        ) 
    ;
    `r[3*10-1:0] SIN_ADRs_Ds     ;
    `ack
        `xar
                                    SIN_ADRs_Ds <= 0 ;
        else
            if( CK_EE_i )           SIN_ADRs_Ds <= {SIN_ADRs_Ds ,sin_adr_s} ;
    `w`s[12:0] sin_dat_s = SIN_ROM_DATs + {SIN_ADRs_Ds[2*10+:10] , 1'b0} ;

    `r[ 2:0]    MINUS_Ds    ;
    `r[ 2:0]    MAX_MIN_Ds  ;
    `r[ 2:0]    ZERO_Ds     ;
    `r`s[11:0]  SINs        ;
    `w[7:0] B_ROM_DLYs = B_ROM_DAT_DLYs - B_IN_DAT_DLYs_i ;
    `r          SIN_CODE_DONE_D ;
    `ack
        `xar
        `b
                                    SINs <= 0 ;
                                    SIN_CODE_DONE_D <= 1'b0 ;
        `eelse 
        `b
                                    SIN_CODE_DONE_D <= SIN_CODE_DONE ;
             if( SIN_CODE_DONE  )
            `b
                if( ZERO_Ds[B_ROM_DLYs-1] )
                                    SINs <= 12'd0 ;
                else
                `b  if(MAX_MIN_Ds[B_ROM_DLYs-1] | (|sin_dat_s[12:11]))
                    `b  if( MINUS_Ds[B_ROM_DLYs-1])
                                    SINs <= -12'h7FF ;
                        else
                                    SINs <=  12'h7FF ;
                    `e else if( MINUS_Ds[B_ROM_DLYs-1] )
                                    SINs <= -sin_dat_s ;
                    else
                                    SINs <=  sin_dat_s ;
                `e
            `e
        `e
    `a SINs_o = SINs ;
    `a DONE_o = SIN_CODE_DONE_D ;
    // ctl
    `ack
        `xar
        `b  MINUS_Ds    <= 0 ;
            MAX_MIN_Ds  <= 0 ;
            ZERO_Ds     <= 1'b1 ;
        `e else if( CK_EE_i )
        `b  MINUS_Ds    <= {MINUS_Ds   ,  DATs_i[11]} ;
            MAX_MIN_Ds  <= {MAX_MIN_Ds , (DATs_i[9:0] == 'd0)} ;
            ZERO_Ds     <= {ZERO_Ds    , (DATs_i[10:0] == 'd0) } ;
        `e
    `a B_OUT_DAT_DLYs_o = B_ROM_DAT_DLYs + C_DAT_DLYs ;
endmodule // SIN_S11_S11
`define SIN_S11_S11
`endif

`ifndef SIN_ROM_S11_S11
// 2ck dly
module SIN_ROM_S11_S11
(     `in`tri1          CK_i
    , `in`tri1          XARST_i
    , `in`tri1          CK_EE_i
    , `in`tri0[7:0]     B_IN_DAT_DLYs_i
    , `in`tri0[ 9:0]    ADRs_i
    , `out`w  [ 8:0]    QQs_o
    , `out`w            DONE_o
    , `out`w[7:0]       B_OUT_DAT_DLYs_o
) ;
    localparam C_DAT_DLYs = 3 ;
    `r [ 9:0]ROM_ADRs ;
    `r  CK_EE_D ;
    `ack
        `xar
        `b
            ROM_ADRs <= 0 ;
            CK_EE_D <= 1'b0 ;
        `eelse 
        `b
            CK_EE_D <= CK_EE_i ;
            if( CK_EE_i )
                ROM_ADRs <= ADRs_i ;
        `e
    // sin_tb_12_12_inc.v
    // datetime.datetime(2015, 12, 20, 11, 29, 28, 266222)
    `r[ 8:0]    QQs ;
    `r          CK_EE_DD ;
    `ack
        `xar
        `b
            QQs <= 0 ;
            CK_EE_DD <= 1'b0 ;
        `eelse
        `b 
            CK_EE_DD <= CK_EE_D ;
            if( CK_EE_D )
            case ( ROM_ADRs )
                10'h000 : QQs <= 9'h000 ;
                10'h001 : QQs <= 9'h001 ;
                10'h002 : QQs <= 9'h002 ;
                10'h003 : QQs <= 9'h003 ;
                10'h004 : QQs <= 9'h005 ;
                10'h005 : QQs <= 9'h006 ;
                10'h006 : QQs <= 9'h007 ;
                10'h007 : QQs <= 9'h008 ;
                10'h008 : QQs <= 9'h009 ;
                10'h009 : QQs <= 9'h00A ;
                10'h00A : QQs <= 9'h00B ;
                10'h00B : QQs <= 9'h00D ;
                10'h00C : QQs <= 9'h00E ;
                10'h00D : QQs <= 9'h00F ;
                10'h00E : QQs <= 9'h010 ;
                10'h00F : QQs <= 9'h011 ;
                10'h010 : QQs <= 9'h012 ;
                10'h011 : QQs <= 9'h013 ;
                10'h012 : QQs <= 9'h015 ;
                10'h013 : QQs <= 9'h016 ;
                10'h014 : QQs <= 9'h017 ;
                10'h015 : QQs <= 9'h018 ;
                10'h016 : QQs <= 9'h019 ;
                10'h017 : QQs <= 9'h01A ;
                10'h018 : QQs <= 9'h01B ;
                10'h019 : QQs <= 9'h01D ;
                10'h01A : QQs <= 9'h01E ;
                10'h01B : QQs <= 9'h01F ;
                10'h01C : QQs <= 9'h020 ;
                10'h01D : QQs <= 9'h021 ;
                10'h01E : QQs <= 9'h022 ;
                10'h01F : QQs <= 9'h023 ;
                10'h020 : QQs <= 9'h024 ;
                10'h021 : QQs <= 9'h026 ;
                10'h022 : QQs <= 9'h027 ;
                10'h023 : QQs <= 9'h028 ;
                10'h024 : QQs <= 9'h029 ;
                10'h025 : QQs <= 9'h02A ;
                10'h026 : QQs <= 9'h02B ;
                10'h027 : QQs <= 9'h02C ;
                10'h028 : QQs <= 9'h02E ;
                10'h029 : QQs <= 9'h02F ;
                10'h02A : QQs <= 9'h030 ;
                10'h02B : QQs <= 9'h031 ;
                10'h02C : QQs <= 9'h032 ;
                10'h02D : QQs <= 9'h033 ;
                10'h02E : QQs <= 9'h034 ;
                10'h02F : QQs <= 9'h036 ;
                10'h030 : QQs <= 9'h037 ;
                10'h031 : QQs <= 9'h038 ;
                10'h032 : QQs <= 9'h039 ;
                10'h033 : QQs <= 9'h03A ;
                10'h034 : QQs <= 9'h03B ;
                10'h035 : QQs <= 9'h03C ;
                10'h036 : QQs <= 9'h03D ;
                10'h037 : QQs <= 9'h03F ;
                10'h038 : QQs <= 9'h040 ;
                10'h039 : QQs <= 9'h041 ;
                10'h03A : QQs <= 9'h042 ;
                10'h03B : QQs <= 9'h043 ;
                10'h03C : QQs <= 9'h044 ;
                10'h03D : QQs <= 9'h045 ;
                10'h03E : QQs <= 9'h046 ;
                10'h03F : QQs <= 9'h048 ;
                10'h040 : QQs <= 9'h049 ;
                10'h041 : QQs <= 9'h04A ;
                10'h042 : QQs <= 9'h04B ;
                10'h043 : QQs <= 9'h04C ;
                10'h044 : QQs <= 9'h04D ;
                10'h045 : QQs <= 9'h04E ;
                10'h046 : QQs <= 9'h04F ;
                10'h047 : QQs <= 9'h051 ;
                10'h048 : QQs <= 9'h052 ;
                10'h049 : QQs <= 9'h053 ;
                10'h04A : QQs <= 9'h054 ;
                10'h04B : QQs <= 9'h055 ;
                10'h04C : QQs <= 9'h056 ;
                10'h04D : QQs <= 9'h057 ;
                10'h04E : QQs <= 9'h058 ;
                10'h04F : QQs <= 9'h05A ;
                10'h050 : QQs <= 9'h05B ;
                10'h051 : QQs <= 9'h05C ;
                10'h052 : QQs <= 9'h05D ;
                10'h053 : QQs <= 9'h05E ;
                10'h054 : QQs <= 9'h05F ;
                10'h055 : QQs <= 9'h060 ;
                10'h056 : QQs <= 9'h061 ;
                10'h057 : QQs <= 9'h063 ;
                10'h058 : QQs <= 9'h064 ;
                10'h059 : QQs <= 9'h065 ;
                10'h05A : QQs <= 9'h066 ;
                10'h05B : QQs <= 9'h067 ;
                10'h05C : QQs <= 9'h068 ;
                10'h05D : QQs <= 9'h069 ;
                10'h05E : QQs <= 9'h06A ;
                10'h05F : QQs <= 9'h06B ;
                10'h060 : QQs <= 9'h06D ;
                10'h061 : QQs <= 9'h06E ;
                10'h062 : QQs <= 9'h06F ;
                10'h063 : QQs <= 9'h070 ;
                10'h064 : QQs <= 9'h071 ;
                10'h065 : QQs <= 9'h072 ;
                10'h066 : QQs <= 9'h073 ;
                10'h067 : QQs <= 9'h074 ;
                10'h068 : QQs <= 9'h075 ;
                10'h069 : QQs <= 9'h076 ;
                10'h06A : QQs <= 9'h078 ;
                10'h06B : QQs <= 9'h079 ;
                10'h06C : QQs <= 9'h07A ;
                10'h06D : QQs <= 9'h07B ;
                10'h06E : QQs <= 9'h07C ;
                10'h06F : QQs <= 9'h07D ;
                10'h070 : QQs <= 9'h07E ;
                10'h071 : QQs <= 9'h07F ;
                10'h072 : QQs <= 9'h080 ;
                10'h073 : QQs <= 9'h081 ;
                10'h074 : QQs <= 9'h083 ;
                10'h075 : QQs <= 9'h084 ;
                10'h076 : QQs <= 9'h085 ;
                10'h077 : QQs <= 9'h086 ;
                10'h078 : QQs <= 9'h087 ;
                10'h079 : QQs <= 9'h088 ;
                10'h07A : QQs <= 9'h089 ;
                10'h07B : QQs <= 9'h08A ;
                10'h07C : QQs <= 9'h08B ;
                10'h07D : QQs <= 9'h08C ;
                10'h07E : QQs <= 9'h08D ;
                10'h07F : QQs <= 9'h08E ;
                10'h080 : QQs <= 9'h090 ;
                10'h081 : QQs <= 9'h091 ;
                10'h082 : QQs <= 9'h092 ;
                10'h083 : QQs <= 9'h093 ;
                10'h084 : QQs <= 9'h094 ;
                10'h085 : QQs <= 9'h095 ;
                10'h086 : QQs <= 9'h096 ;
                10'h087 : QQs <= 9'h097 ;
                10'h088 : QQs <= 9'h098 ;
                10'h089 : QQs <= 9'h099 ;
                10'h08A : QQs <= 9'h09A ;
                10'h08B : QQs <= 9'h09B ;
                10'h08C : QQs <= 9'h09C ;
                10'h08D : QQs <= 9'h09E ;
                10'h08E : QQs <= 9'h09F ;
                10'h08F : QQs <= 9'h0A0 ;
                10'h090 : QQs <= 9'h0A1 ;
                10'h091 : QQs <= 9'h0A2 ;
                10'h092 : QQs <= 9'h0A3 ;
                10'h093 : QQs <= 9'h0A4 ;
                10'h094 : QQs <= 9'h0A5 ;
                10'h095 : QQs <= 9'h0A6 ;
                10'h096 : QQs <= 9'h0A7 ;
                10'h097 : QQs <= 9'h0A8 ;
                10'h098 : QQs <= 9'h0A9 ;
                10'h099 : QQs <= 9'h0AA ;
                10'h09A : QQs <= 9'h0AB ;
                10'h09B : QQs <= 9'h0AC ;
                10'h09C : QQs <= 9'h0AD ;
                10'h09D : QQs <= 9'h0AE ;
                10'h09E : QQs <= 9'h0B0 ;
                10'h09F : QQs <= 9'h0B1 ;
                10'h0A0 : QQs <= 9'h0B2 ;
                10'h0A1 : QQs <= 9'h0B3 ;
                10'h0A2 : QQs <= 9'h0B4 ;
                10'h0A3 : QQs <= 9'h0B5 ;
                10'h0A4 : QQs <= 9'h0B6 ;
                10'h0A5 : QQs <= 9'h0B7 ;
                10'h0A6 : QQs <= 9'h0B8 ;
                10'h0A7 : QQs <= 9'h0B9 ;
                10'h0A8 : QQs <= 9'h0BA ;
                10'h0A9 : QQs <= 9'h0BB ;
                10'h0AA : QQs <= 9'h0BC ;
                10'h0AB : QQs <= 9'h0BD ;
                10'h0AC : QQs <= 9'h0BE ;
                10'h0AD : QQs <= 9'h0BF ;
                10'h0AE : QQs <= 9'h0C0 ;
                10'h0AF : QQs <= 9'h0C1 ;
                10'h0B0 : QQs <= 9'h0C2 ;
                10'h0B1 : QQs <= 9'h0C3 ;
                10'h0B2 : QQs <= 9'h0C4 ;
                10'h0B3 : QQs <= 9'h0C5 ;
                10'h0B4 : QQs <= 9'h0C6 ;
                10'h0B5 : QQs <= 9'h0C7 ;
                10'h0B6 : QQs <= 9'h0C8 ;
                10'h0B7 : QQs <= 9'h0C9 ;
                10'h0B8 : QQs <= 9'h0CA ;
                10'h0B9 : QQs <= 9'h0CB ;
                10'h0BA : QQs <= 9'h0CC ;
                10'h0BB : QQs <= 9'h0CD ;
                10'h0BC : QQs <= 9'h0CE ;
                10'h0BD : QQs <= 9'h0CF ;
                10'h0BE : QQs <= 9'h0D0 ;
                10'h0BF : QQs <= 9'h0D1 ;
                10'h0C0 : QQs <= 9'h0D3 ;
                10'h0C1 : QQs <= 9'h0D4 ;
                10'h0C2 : QQs <= 9'h0D5 ;
                10'h0C3 : QQs <= 9'h0D6 ;
                10'h0C4 : QQs <= 9'h0D7 ;
                10'h0C5 : QQs <= 9'h0D8 ;
                10'h0C6 : QQs <= 9'h0D9 ;
                10'h0C7 : QQs <= 9'h0DA ;
                10'h0C8 : QQs <= 9'h0DB ;
                10'h0C9 : QQs <= 9'h0DC ;
                10'h0CA : QQs <= 9'h0DC ;
                10'h0CB : QQs <= 9'h0DD ;
                10'h0CC : QQs <= 9'h0DE ;
                10'h0CD : QQs <= 9'h0DF ;
                10'h0CE : QQs <= 9'h0E0 ;
                10'h0CF : QQs <= 9'h0E1 ;
                10'h0D0 : QQs <= 9'h0E2 ;
                10'h0D1 : QQs <= 9'h0E3 ;
                10'h0D2 : QQs <= 9'h0E4 ;
                10'h0D3 : QQs <= 9'h0E5 ;
                10'h0D4 : QQs <= 9'h0E6 ;
                10'h0D5 : QQs <= 9'h0E7 ;
                10'h0D6 : QQs <= 9'h0E8 ;
                10'h0D7 : QQs <= 9'h0E9 ;
                10'h0D8 : QQs <= 9'h0EA ;
                10'h0D9 : QQs <= 9'h0EB ;
                10'h0DA : QQs <= 9'h0EC ;
                10'h0DB : QQs <= 9'h0ED ;
                10'h0DC : QQs <= 9'h0EE ;
                10'h0DD : QQs <= 9'h0EF ;
                10'h0DE : QQs <= 9'h0F0 ;
                10'h0DF : QQs <= 9'h0F1 ;
                10'h0E0 : QQs <= 9'h0F2 ;
                10'h0E1 : QQs <= 9'h0F3 ;
                10'h0E2 : QQs <= 9'h0F4 ;
                10'h0E3 : QQs <= 9'h0F5 ;
                10'h0E4 : QQs <= 9'h0F6 ;
                10'h0E5 : QQs <= 9'h0F7 ;
                10'h0E6 : QQs <= 9'h0F8 ;
                10'h0E7 : QQs <= 9'h0F9 ;
                10'h0E8 : QQs <= 9'h0FA ;
                10'h0E9 : QQs <= 9'h0FB ;
                10'h0EA : QQs <= 9'h0FB ;
                10'h0EB : QQs <= 9'h0FC ;
                10'h0EC : QQs <= 9'h0FD ;
                10'h0ED : QQs <= 9'h0FE ;
                10'h0EE : QQs <= 9'h0FF ;
                10'h0EF : QQs <= 9'h100 ;
                10'h0F0 : QQs <= 9'h101 ;
                10'h0F1 : QQs <= 9'h102 ;
                10'h0F2 : QQs <= 9'h103 ;
                10'h0F3 : QQs <= 9'h104 ;
                10'h0F4 : QQs <= 9'h105 ;
                10'h0F5 : QQs <= 9'h106 ;
                10'h0F6 : QQs <= 9'h107 ;
                10'h0F7 : QQs <= 9'h108 ;
                10'h0F8 : QQs <= 9'h108 ;
                10'h0F9 : QQs <= 9'h109 ;
                10'h0FA : QQs <= 9'h10A ;
                10'h0FB : QQs <= 9'h10B ;
                10'h0FC : QQs <= 9'h10C ;
                10'h0FD : QQs <= 9'h10D ;
                10'h0FE : QQs <= 9'h10E ;
                10'h0FF : QQs <= 9'h10F ;
                10'h100 : QQs <= 9'h110 ;
                10'h101 : QQs <= 9'h111 ;
                10'h102 : QQs <= 9'h112 ;
                10'h103 : QQs <= 9'h112 ;
                10'h104 : QQs <= 9'h113 ;
                10'h105 : QQs <= 9'h114 ;
                10'h106 : QQs <= 9'h115 ;
                10'h107 : QQs <= 9'h116 ;
                10'h108 : QQs <= 9'h117 ;
                10'h109 : QQs <= 9'h118 ;
                10'h10A : QQs <= 9'h119 ;
                10'h10B : QQs <= 9'h11A ;
                10'h10C : QQs <= 9'h11A ;
                10'h10D : QQs <= 9'h11B ;
                10'h10E : QQs <= 9'h11C ;
                10'h10F : QQs <= 9'h11D ;
                10'h110 : QQs <= 9'h11E ;
                10'h111 : QQs <= 9'h11F ;
                10'h112 : QQs <= 9'h120 ;
                10'h113 : QQs <= 9'h121 ;
                10'h114 : QQs <= 9'h121 ;
                10'h115 : QQs <= 9'h122 ;
                10'h116 : QQs <= 9'h123 ;
                10'h117 : QQs <= 9'h124 ;
                10'h118 : QQs <= 9'h125 ;
                10'h119 : QQs <= 9'h126 ;
                10'h11A : QQs <= 9'h127 ;
                10'h11B : QQs <= 9'h127 ;
                10'h11C : QQs <= 9'h128 ;
                10'h11D : QQs <= 9'h129 ;
                10'h11E : QQs <= 9'h12A ;
                10'h11F : QQs <= 9'h12B ;
                10'h120 : QQs <= 9'h12C ;
                10'h121 : QQs <= 9'h12C ;
                10'h122 : QQs <= 9'h12D ;
                10'h123 : QQs <= 9'h12E ;
                10'h124 : QQs <= 9'h12F ;
                10'h125 : QQs <= 9'h130 ;
                10'h126 : QQs <= 9'h131 ;
                10'h127 : QQs <= 9'h131 ;
                10'h128 : QQs <= 9'h132 ;
                10'h129 : QQs <= 9'h133 ;
                10'h12A : QQs <= 9'h134 ;
                10'h12B : QQs <= 9'h135 ;
                10'h12C : QQs <= 9'h136 ;
                10'h12D : QQs <= 9'h136 ;
                10'h12E : QQs <= 9'h137 ;
                10'h12F : QQs <= 9'h138 ;
                10'h130 : QQs <= 9'h139 ;
                10'h131 : QQs <= 9'h13A ;
                10'h132 : QQs <= 9'h13A ;
                10'h133 : QQs <= 9'h13B ;
                10'h134 : QQs <= 9'h13C ;
                10'h135 : QQs <= 9'h13D ;
                10'h136 : QQs <= 9'h13E ;
                10'h137 : QQs <= 9'h13E ;
                10'h138 : QQs <= 9'h13F ;
                10'h139 : QQs <= 9'h140 ;
                10'h13A : QQs <= 9'h141 ;
                10'h13B : QQs <= 9'h142 ;
                10'h13C : QQs <= 9'h142 ;
                10'h13D : QQs <= 9'h143 ;
                10'h13E : QQs <= 9'h144 ;
                10'h13F : QQs <= 9'h145 ;
                10'h140 : QQs <= 9'h145 ;
                10'h141 : QQs <= 9'h146 ;
                10'h142 : QQs <= 9'h147 ;
                10'h143 : QQs <= 9'h148 ;
                10'h144 : QQs <= 9'h148 ;
                10'h145 : QQs <= 9'h149 ;
                10'h146 : QQs <= 9'h14A ;
                10'h147 : QQs <= 9'h14B ;
                10'h148 : QQs <= 9'h14C ;
                10'h149 : QQs <= 9'h14C ;
                10'h14A : QQs <= 9'h14D ;
                10'h14B : QQs <= 9'h14E ;
                10'h14C : QQs <= 9'h14F ;
                10'h14D : QQs <= 9'h14F ;
                10'h14E : QQs <= 9'h150 ;
                10'h14F : QQs <= 9'h151 ;
                10'h150 : QQs <= 9'h151 ;
                10'h151 : QQs <= 9'h152 ;
                10'h152 : QQs <= 9'h153 ;
                10'h153 : QQs <= 9'h154 ;
                10'h154 : QQs <= 9'h154 ;
                10'h155 : QQs <= 9'h155 ;
                10'h156 : QQs <= 9'h156 ;
                10'h157 : QQs <= 9'h157 ;
                10'h158 : QQs <= 9'h157 ;
                10'h159 : QQs <= 9'h158 ;
                10'h15A : QQs <= 9'h159 ;
                10'h15B : QQs <= 9'h159 ;
                10'h15C : QQs <= 9'h15A ;
                10'h15D : QQs <= 9'h15B ;
                10'h15E : QQs <= 9'h15B ;
                10'h15F : QQs <= 9'h15C ;
                10'h160 : QQs <= 9'h15D ;
                10'h161 : QQs <= 9'h15E ;
                10'h162 : QQs <= 9'h15E ;
                10'h163 : QQs <= 9'h15F ;
                10'h164 : QQs <= 9'h160 ;
                10'h165 : QQs <= 9'h160 ;
                10'h166 : QQs <= 9'h161 ;
                10'h167 : QQs <= 9'h162 ;
                10'h168 : QQs <= 9'h162 ;
                10'h169 : QQs <= 9'h163 ;
                10'h16A : QQs <= 9'h164 ;
                10'h16B : QQs <= 9'h164 ;
                10'h16C : QQs <= 9'h165 ;
                10'h16D : QQs <= 9'h166 ;
                10'h16E : QQs <= 9'h166 ;
                10'h16F : QQs <= 9'h167 ;
                10'h170 : QQs <= 9'h168 ;
                10'h171 : QQs <= 9'h168 ;
                10'h172 : QQs <= 9'h169 ;
                10'h173 : QQs <= 9'h16A ;
                10'h174 : QQs <= 9'h16A ;
                10'h175 : QQs <= 9'h16B ;
                10'h176 : QQs <= 9'h16C ;
                10'h177 : QQs <= 9'h16C ;
                10'h178 : QQs <= 9'h16D ;
                10'h179 : QQs <= 9'h16D ;
                10'h17A : QQs <= 9'h16E ;
                10'h17B : QQs <= 9'h16F ;
                10'h17C : QQs <= 9'h16F ;
                10'h17D : QQs <= 9'h170 ;
                10'h17E : QQs <= 9'h171 ;
                10'h17F : QQs <= 9'h171 ;
                10'h180 : QQs <= 9'h172 ;
                10'h181 : QQs <= 9'h172 ;
                10'h182 : QQs <= 9'h173 ;
                10'h183 : QQs <= 9'h174 ;
                10'h184 : QQs <= 9'h174 ;
                10'h185 : QQs <= 9'h175 ;
                10'h186 : QQs <= 9'h175 ;
                10'h187 : QQs <= 9'h176 ;
                10'h188 : QQs <= 9'h177 ;
                10'h189 : QQs <= 9'h177 ;
                10'h18A : QQs <= 9'h178 ;
                10'h18B : QQs <= 9'h178 ;
                10'h18C : QQs <= 9'h179 ;
                10'h18D : QQs <= 9'h17A ;
                10'h18E : QQs <= 9'h17A ;
                10'h18F : QQs <= 9'h17B ;
                10'h190 : QQs <= 9'h17B ;
                10'h191 : QQs <= 9'h17C ;
                10'h192 : QQs <= 9'h17C ;
                10'h193 : QQs <= 9'h17D ;
                10'h194 : QQs <= 9'h17E ;
                10'h195 : QQs <= 9'h17E ;
                10'h196 : QQs <= 9'h17F ;
                10'h197 : QQs <= 9'h17F ;
                10'h198 : QQs <= 9'h180 ;
                10'h199 : QQs <= 9'h180 ;
                10'h19A : QQs <= 9'h181 ;
                10'h19B : QQs <= 9'h181 ;
                10'h19C : QQs <= 9'h182 ;
                10'h19D : QQs <= 9'h182 ;
                10'h19E : QQs <= 9'h183 ;
                10'h19F : QQs <= 9'h183 ;
                10'h1A0 : QQs <= 9'h184 ;
                10'h1A1 : QQs <= 9'h185 ;
                10'h1A2 : QQs <= 9'h185 ;
                10'h1A3 : QQs <= 9'h186 ;
                10'h1A4 : QQs <= 9'h186 ;
                10'h1A5 : QQs <= 9'h187 ;
                10'h1A6 : QQs <= 9'h187 ;
                10'h1A7 : QQs <= 9'h188 ;
                10'h1A8 : QQs <= 9'h188 ;
                10'h1A9 : QQs <= 9'h189 ;
                10'h1AA : QQs <= 9'h189 ;
                10'h1AB : QQs <= 9'h18A ;
                10'h1AC : QQs <= 9'h18A ;
                10'h1AD : QQs <= 9'h18B ;
                10'h1AE : QQs <= 9'h18B ;
                10'h1AF : QQs <= 9'h18C ;
                10'h1B0 : QQs <= 9'h18C ;
                10'h1B1 : QQs <= 9'h18C ;
                10'h1B2 : QQs <= 9'h18D ;
                10'h1B3 : QQs <= 9'h18D ;
                10'h1B4 : QQs <= 9'h18E ;
                10'h1B5 : QQs <= 9'h18E ;
                10'h1B6 : QQs <= 9'h18F ;
                10'h1B7 : QQs <= 9'h18F ;
                10'h1B8 : QQs <= 9'h190 ;
                10'h1B9 : QQs <= 9'h190 ;
                10'h1BA : QQs <= 9'h191 ;
                10'h1BB : QQs <= 9'h191 ;
                10'h1BC : QQs <= 9'h191 ;
                10'h1BD : QQs <= 9'h192 ;
                10'h1BE : QQs <= 9'h192 ;
                10'h1BF : QQs <= 9'h193 ;
                10'h1C0 : QQs <= 9'h193 ;
                10'h1C1 : QQs <= 9'h194 ;
                10'h1C2 : QQs <= 9'h194 ;
                10'h1C3 : QQs <= 9'h195 ;
                10'h1C4 : QQs <= 9'h195 ;
                10'h1C5 : QQs <= 9'h195 ;
                10'h1C6 : QQs <= 9'h196 ;
                10'h1C7 : QQs <= 9'h196 ;
                10'h1C8 : QQs <= 9'h197 ;
                10'h1C9 : QQs <= 9'h197 ;
                10'h1CA : QQs <= 9'h197 ;
                10'h1CB : QQs <= 9'h198 ;
                10'h1CC : QQs <= 9'h198 ;
                10'h1CD : QQs <= 9'h199 ;
                10'h1CE : QQs <= 9'h199 ;
                10'h1CF : QQs <= 9'h199 ;
                10'h1D0 : QQs <= 9'h19A ;
                10'h1D1 : QQs <= 9'h19A ;
                10'h1D2 : QQs <= 9'h19A ;
                10'h1D3 : QQs <= 9'h19B ;
                10'h1D4 : QQs <= 9'h19B ;
                10'h1D5 : QQs <= 9'h19C ;
                10'h1D6 : QQs <= 9'h19C ;
                10'h1D7 : QQs <= 9'h19C ;
                10'h1D8 : QQs <= 9'h19D ;
                10'h1D9 : QQs <= 9'h19D ;
                10'h1DA : QQs <= 9'h19D ;
                10'h1DB : QQs <= 9'h19E ;
                10'h1DC : QQs <= 9'h19E ;
                10'h1DD : QQs <= 9'h19E ;
                10'h1DE : QQs <= 9'h19F ;
                10'h1DF : QQs <= 9'h19F ;
                10'h1E0 : QQs <= 9'h19F ;
                10'h1E1 : QQs <= 9'h1A0 ;
                10'h1E2 : QQs <= 9'h1A0 ;
                10'h1E3 : QQs <= 9'h1A0 ;
                10'h1E4 : QQs <= 9'h1A1 ;
                10'h1E5 : QQs <= 9'h1A1 ;
                10'h1E6 : QQs <= 9'h1A1 ;
                10'h1E7 : QQs <= 9'h1A2 ;
                10'h1E8 : QQs <= 9'h1A2 ;
                10'h1E9 : QQs <= 9'h1A2 ;
                10'h1EA : QQs <= 9'h1A2 ;
                10'h1EB : QQs <= 9'h1A3 ;
                10'h1EC : QQs <= 9'h1A3 ;
                10'h1ED : QQs <= 9'h1A3 ;
                10'h1EE : QQs <= 9'h1A4 ;
                10'h1EF : QQs <= 9'h1A4 ;
                10'h1F0 : QQs <= 9'h1A4 ;
                10'h1F1 : QQs <= 9'h1A4 ;
                10'h1F2 : QQs <= 9'h1A5 ;
                10'h1F3 : QQs <= 9'h1A5 ;
                10'h1F4 : QQs <= 9'h1A5 ;
                10'h1F5 : QQs <= 9'h1A6 ;
                10'h1F6 : QQs <= 9'h1A6 ;
                10'h1F7 : QQs <= 9'h1A6 ;
                10'h1F8 : QQs <= 9'h1A6 ;
                10'h1F9 : QQs <= 9'h1A7 ;
                10'h1FA : QQs <= 9'h1A7 ;
                10'h1FB : QQs <= 9'h1A7 ;
                10'h1FC : QQs <= 9'h1A7 ;
                10'h1FD : QQs <= 9'h1A7 ;
                10'h1FE : QQs <= 9'h1A8 ;
                10'h1FF : QQs <= 9'h1A8 ;
                10'h200 : QQs <= 9'h1A8 ;
                10'h201 : QQs <= 9'h1A8 ;
                10'h202 : QQs <= 9'h1A9 ;
                10'h203 : QQs <= 9'h1A9 ;
                10'h204 : QQs <= 9'h1A9 ;
                10'h205 : QQs <= 9'h1A9 ;
                10'h206 : QQs <= 9'h1A9 ;
                10'h207 : QQs <= 9'h1AA ;
                10'h208 : QQs <= 9'h1AA ;
                10'h209 : QQs <= 9'h1AA ;
                10'h20A : QQs <= 9'h1AA ;
                10'h20B : QQs <= 9'h1AA ;
                10'h20C : QQs <= 9'h1AB ;
                10'h20D : QQs <= 9'h1AB ;
                10'h20E : QQs <= 9'h1AB ;
                10'h20F : QQs <= 9'h1AB ;
                10'h210 : QQs <= 9'h1AB ;
                10'h211 : QQs <= 9'h1AB ;
                10'h212 : QQs <= 9'h1AC ;
                10'h213 : QQs <= 9'h1AC ;
                10'h214 : QQs <= 9'h1AC ;
                10'h215 : QQs <= 9'h1AC ;
                10'h216 : QQs <= 9'h1AC ;
                10'h217 : QQs <= 9'h1AC ;
                10'h218 : QQs <= 9'h1AC ;
                10'h219 : QQs <= 9'h1AD ;
                10'h21A : QQs <= 9'h1AD ;
                10'h21B : QQs <= 9'h1AD ;
                10'h21C : QQs <= 9'h1AD ;
                10'h21D : QQs <= 9'h1AD ;
                10'h21E : QQs <= 9'h1AD ;
                10'h21F : QQs <= 9'h1AD ;
                10'h220 : QQs <= 9'h1AD ;
                10'h221 : QQs <= 9'h1AE ;
                10'h222 : QQs <= 9'h1AE ;
                10'h223 : QQs <= 9'h1AE ;
                10'h224 : QQs <= 9'h1AE ;
                10'h225 : QQs <= 9'h1AE ;
                10'h226 : QQs <= 9'h1AE ;
                10'h227 : QQs <= 9'h1AE ;
                10'h228 : QQs <= 9'h1AE ;
                10'h229 : QQs <= 9'h1AE ;
                10'h22A : QQs <= 9'h1AE ;
                10'h22B : QQs <= 9'h1AE ;
                10'h22C : QQs <= 9'h1AF ;
                10'h22D : QQs <= 9'h1AF ;
                10'h22E : QQs <= 9'h1AF ;
                10'h22F : QQs <= 9'h1AF ;
                10'h230 : QQs <= 9'h1AF ;
                10'h231 : QQs <= 9'h1AF ;
                10'h232 : QQs <= 9'h1AF ;
                10'h233 : QQs <= 9'h1AF ;
                10'h234 : QQs <= 9'h1AF ;
                10'h235 : QQs <= 9'h1AF ;
                10'h236 : QQs <= 9'h1AF ;
                10'h237 : QQs <= 9'h1AF ;
                10'h238 : QQs <= 9'h1AF ;
                10'h239 : QQs <= 9'h1AF ;
                10'h23A : QQs <= 9'h1AF ;
                10'h23B : QQs <= 9'h1AF ;
                10'h23C : QQs <= 9'h1AF ;
                10'h23D : QQs <= 9'h1AF ;
                10'h23E : QQs <= 9'h1AF ;
                10'h23F : QQs <= 9'h1AF ;
                10'h240 : QQs <= 9'h1AF ;
                10'h241 : QQs <= 9'h1AF ;
                10'h242 : QQs <= 9'h1AF ;
                10'h243 : QQs <= 9'h1AF ;
                10'h244 : QQs <= 9'h1AF ;
                10'h245 : QQs <= 9'h1AF ;
                10'h246 : QQs <= 9'h1AF ;
                10'h247 : QQs <= 9'h1AF ;
                10'h248 : QQs <= 9'h1AF ;
                10'h249 : QQs <= 9'h1AF ;
                10'h24A : QQs <= 9'h1AF ;
                10'h24B : QQs <= 9'h1AF ;
                10'h24C : QQs <= 9'h1AF ;
                10'h24D : QQs <= 9'h1AF ;
                10'h24E : QQs <= 9'h1AF ;
                10'h24F : QQs <= 9'h1AF ;
                10'h250 : QQs <= 9'h1AF ;
                10'h251 : QQs <= 9'h1AE ;
                10'h252 : QQs <= 9'h1AE ;
                10'h253 : QQs <= 9'h1AE ;
                10'h254 : QQs <= 9'h1AE ;
                10'h255 : QQs <= 9'h1AE ;
                10'h256 : QQs <= 9'h1AE ;
                10'h257 : QQs <= 9'h1AE ;
                10'h258 : QQs <= 9'h1AE ;
                10'h259 : QQs <= 9'h1AE ;
                10'h25A : QQs <= 9'h1AE ;
                10'h25B : QQs <= 9'h1AE ;
                10'h25C : QQs <= 9'h1AD ;
                10'h25D : QQs <= 9'h1AD ;
                10'h25E : QQs <= 9'h1AD ;
                10'h25F : QQs <= 9'h1AD ;
                10'h260 : QQs <= 9'h1AD ;
                10'h261 : QQs <= 9'h1AD ;
                10'h262 : QQs <= 9'h1AD ;
                10'h263 : QQs <= 9'h1AD ;
                10'h264 : QQs <= 9'h1AC ;
                10'h265 : QQs <= 9'h1AC ;
                10'h266 : QQs <= 9'h1AC ;
                10'h267 : QQs <= 9'h1AC ;
                10'h268 : QQs <= 9'h1AC ;
                10'h269 : QQs <= 9'h1AC ;
                10'h26A : QQs <= 9'h1AB ;
                10'h26B : QQs <= 9'h1AB ;
                10'h26C : QQs <= 9'h1AB ;
                10'h26D : QQs <= 9'h1AB ;
                10'h26E : QQs <= 9'h1AB ;
                10'h26F : QQs <= 9'h1AB ;
                10'h270 : QQs <= 9'h1AA ;
                10'h271 : QQs <= 9'h1AA ;
                10'h272 : QQs <= 9'h1AA ;
                10'h273 : QQs <= 9'h1AA ;
                10'h274 : QQs <= 9'h1AA ;
                10'h275 : QQs <= 9'h1A9 ;
                10'h276 : QQs <= 9'h1A9 ;
                10'h277 : QQs <= 9'h1A9 ;
                10'h278 : QQs <= 9'h1A9 ;
                10'h279 : QQs <= 9'h1A9 ;
                10'h27A : QQs <= 9'h1A8 ;
                10'h27B : QQs <= 9'h1A8 ;
                10'h27C : QQs <= 9'h1A8 ;
                10'h27D : QQs <= 9'h1A8 ;
                10'h27E : QQs <= 9'h1A7 ;
                10'h27F : QQs <= 9'h1A7 ;
                10'h280 : QQs <= 9'h1A7 ;
                10'h281 : QQs <= 9'h1A7 ;
                10'h282 : QQs <= 9'h1A6 ;
                10'h283 : QQs <= 9'h1A6 ;
                10'h284 : QQs <= 9'h1A6 ;
                10'h285 : QQs <= 9'h1A6 ;
                10'h286 : QQs <= 9'h1A5 ;
                10'h287 : QQs <= 9'h1A5 ;
                10'h288 : QQs <= 9'h1A5 ;
                10'h289 : QQs <= 9'h1A4 ;
                10'h28A : QQs <= 9'h1A4 ;
                10'h28B : QQs <= 9'h1A4 ;
                10'h28C : QQs <= 9'h1A4 ;
                10'h28D : QQs <= 9'h1A3 ;
                10'h28E : QQs <= 9'h1A3 ;
                10'h28F : QQs <= 9'h1A3 ;
                10'h290 : QQs <= 9'h1A2 ;
                10'h291 : QQs <= 9'h1A2 ;
                10'h292 : QQs <= 9'h1A2 ;
                10'h293 : QQs <= 9'h1A1 ;
                10'h294 : QQs <= 9'h1A1 ;
                10'h295 : QQs <= 9'h1A1 ;
                10'h296 : QQs <= 9'h1A0 ;
                10'h297 : QQs <= 9'h1A0 ;
                10'h298 : QQs <= 9'h1A0 ;
                10'h299 : QQs <= 9'h19F ;
                10'h29A : QQs <= 9'h19F ;
                10'h29B : QQs <= 9'h19F ;
                10'h29C : QQs <= 9'h19E ;
                10'h29D : QQs <= 9'h19E ;
                10'h29E : QQs <= 9'h19D ;
                10'h29F : QQs <= 9'h19D ;
                10'h2A0 : QQs <= 9'h19D ;
                10'h2A1 : QQs <= 9'h19C ;
                10'h2A2 : QQs <= 9'h19C ;
                10'h2A3 : QQs <= 9'h19B ;
                10'h2A4 : QQs <= 9'h19B ;
                10'h2A5 : QQs <= 9'h19B ;
                10'h2A6 : QQs <= 9'h19A ;
                10'h2A7 : QQs <= 9'h19A ;
                10'h2A8 : QQs <= 9'h199 ;
                10'h2A9 : QQs <= 9'h199 ;
                10'h2AA : QQs <= 9'h199 ;
                10'h2AB : QQs <= 9'h198 ;
                10'h2AC : QQs <= 9'h198 ;
                10'h2AD : QQs <= 9'h197 ;
                10'h2AE : QQs <= 9'h197 ;
                10'h2AF : QQs <= 9'h196 ;
                10'h2B0 : QQs <= 9'h196 ;
                10'h2B1 : QQs <= 9'h195 ;
                10'h2B2 : QQs <= 9'h195 ;
                10'h2B3 : QQs <= 9'h195 ;
                10'h2B4 : QQs <= 9'h194 ;
                10'h2B5 : QQs <= 9'h194 ;
                10'h2B6 : QQs <= 9'h193 ;
                10'h2B7 : QQs <= 9'h193 ;
                10'h2B8 : QQs <= 9'h192 ;
                10'h2B9 : QQs <= 9'h192 ;
                10'h2BA : QQs <= 9'h191 ;
                10'h2BB : QQs <= 9'h191 ;
                10'h2BC : QQs <= 9'h190 ;
                10'h2BD : QQs <= 9'h190 ;
                10'h2BE : QQs <= 9'h18F ;
                10'h2BF : QQs <= 9'h18F ;
                10'h2C0 : QQs <= 9'h18E ;
                10'h2C1 : QQs <= 9'h18E ;
                10'h2C2 : QQs <= 9'h18D ;
                10'h2C3 : QQs <= 9'h18D ;
                10'h2C4 : QQs <= 9'h18C ;
                10'h2C5 : QQs <= 9'h18C ;
                10'h2C6 : QQs <= 9'h18B ;
                10'h2C7 : QQs <= 9'h18A ;
                10'h2C8 : QQs <= 9'h18A ;
                10'h2C9 : QQs <= 9'h189 ;
                10'h2CA : QQs <= 9'h189 ;
                10'h2CB : QQs <= 9'h188 ;
                10'h2CC : QQs <= 9'h188 ;
                10'h2CD : QQs <= 9'h187 ;
                10'h2CE : QQs <= 9'h186 ;
                10'h2CF : QQs <= 9'h186 ;
                10'h2D0 : QQs <= 9'h185 ;
                10'h2D1 : QQs <= 9'h185 ;
                10'h2D2 : QQs <= 9'h184 ;
                10'h2D3 : QQs <= 9'h184 ;
                10'h2D4 : QQs <= 9'h183 ;
                10'h2D5 : QQs <= 9'h182 ;
                10'h2D6 : QQs <= 9'h182 ;
                10'h2D7 : QQs <= 9'h181 ;
                10'h2D8 : QQs <= 9'h180 ;
                10'h2D9 : QQs <= 9'h180 ;
                10'h2DA : QQs <= 9'h17F ;
                10'h2DB : QQs <= 9'h17F ;
                10'h2DC : QQs <= 9'h17E ;
                10'h2DD : QQs <= 9'h17D ;
                10'h2DE : QQs <= 9'h17D ;
                10'h2DF : QQs <= 9'h17C ;
                10'h2E0 : QQs <= 9'h17B ;
                10'h2E1 : QQs <= 9'h17B ;
                10'h2E2 : QQs <= 9'h17A ;
                10'h2E3 : QQs <= 9'h179 ;
                10'h2E4 : QQs <= 9'h179 ;
                10'h2E5 : QQs <= 9'h178 ;
                10'h2E6 : QQs <= 9'h177 ;
                10'h2E7 : QQs <= 9'h177 ;
                10'h2E8 : QQs <= 9'h176 ;
                10'h2E9 : QQs <= 9'h175 ;
                10'h2EA : QQs <= 9'h175 ;
                10'h2EB : QQs <= 9'h174 ;
                10'h2EC : QQs <= 9'h173 ;
                10'h2ED : QQs <= 9'h172 ;
                10'h2EE : QQs <= 9'h172 ;
                10'h2EF : QQs <= 9'h171 ;
                10'h2F0 : QQs <= 9'h170 ;
                10'h2F1 : QQs <= 9'h170 ;
                10'h2F2 : QQs <= 9'h16F ;
                10'h2F3 : QQs <= 9'h16E ;
                10'h2F4 : QQs <= 9'h16D ;
                10'h2F5 : QQs <= 9'h16D ;
                10'h2F6 : QQs <= 9'h16C ;
                10'h2F7 : QQs <= 9'h16B ;
                10'h2F8 : QQs <= 9'h16A ;
                10'h2F9 : QQs <= 9'h16A ;
                10'h2FA : QQs <= 9'h169 ;
                10'h2FB : QQs <= 9'h168 ;
                10'h2FC : QQs <= 9'h167 ;
                10'h2FD : QQs <= 9'h166 ;
                10'h2FE : QQs <= 9'h166 ;
                10'h2FF : QQs <= 9'h165 ;
                10'h300 : QQs <= 9'h164 ;
                10'h301 : QQs <= 9'h163 ;
                10'h302 : QQs <= 9'h163 ;
                10'h303 : QQs <= 9'h162 ;
                10'h304 : QQs <= 9'h161 ;
                10'h305 : QQs <= 9'h160 ;
                10'h306 : QQs <= 9'h15F ;
                10'h307 : QQs <= 9'h15E ;
                10'h308 : QQs <= 9'h15E ;
                10'h309 : QQs <= 9'h15D ;
                10'h30A : QQs <= 9'h15C ;
                10'h30B : QQs <= 9'h15B ;
                10'h30C : QQs <= 9'h15A ;
                10'h30D : QQs <= 9'h159 ;
                10'h30E : QQs <= 9'h158 ;
                10'h30F : QQs <= 9'h158 ;
                10'h310 : QQs <= 9'h157 ;
                10'h311 : QQs <= 9'h156 ;
                10'h312 : QQs <= 9'h155 ;
                10'h313 : QQs <= 9'h154 ;
                10'h314 : QQs <= 9'h153 ;
                10'h315 : QQs <= 9'h152 ;
                10'h316 : QQs <= 9'h151 ;
                10'h317 : QQs <= 9'h151 ;
                10'h318 : QQs <= 9'h150 ;
                10'h319 : QQs <= 9'h14F ;
                10'h31A : QQs <= 9'h14E ;
                10'h31B : QQs <= 9'h14D ;
                10'h31C : QQs <= 9'h14C ;
                10'h31D : QQs <= 9'h14B ;
                10'h31E : QQs <= 9'h14A ;
                10'h31F : QQs <= 9'h149 ;
                10'h320 : QQs <= 9'h148 ;
                10'h321 : QQs <= 9'h147 ;
                10'h322 : QQs <= 9'h146 ;
                10'h323 : QQs <= 9'h145 ;
                10'h324 : QQs <= 9'h144 ;
                10'h325 : QQs <= 9'h144 ;
                10'h326 : QQs <= 9'h143 ;
                10'h327 : QQs <= 9'h142 ;
                10'h328 : QQs <= 9'h141 ;
                10'h329 : QQs <= 9'h140 ;
                10'h32A : QQs <= 9'h13F ;
                10'h32B : QQs <= 9'h13E ;
                10'h32C : QQs <= 9'h13D ;
                10'h32D : QQs <= 9'h13C ;
                10'h32E : QQs <= 9'h13B ;
                10'h32F : QQs <= 9'h13A ;
                10'h330 : QQs <= 9'h139 ;
                10'h331 : QQs <= 9'h138 ;
                10'h332 : QQs <= 9'h137 ;
                10'h333 : QQs <= 9'h136 ;
                10'h334 : QQs <= 9'h135 ;
                10'h335 : QQs <= 9'h134 ;
                10'h336 : QQs <= 9'h132 ;
                10'h337 : QQs <= 9'h131 ;
                10'h338 : QQs <= 9'h130 ;
                10'h339 : QQs <= 9'h12F ;
                10'h33A : QQs <= 9'h12E ;
                10'h33B : QQs <= 9'h12D ;
                10'h33C : QQs <= 9'h12C ;
                10'h33D : QQs <= 9'h12B ;
                10'h33E : QQs <= 9'h12A ;
                10'h33F : QQs <= 9'h129 ;
                10'h340 : QQs <= 9'h128 ;
                10'h341 : QQs <= 9'h127 ;
                10'h342 : QQs <= 9'h126 ;
                10'h343 : QQs <= 9'h125 ;
                10'h344 : QQs <= 9'h123 ;
                10'h345 : QQs <= 9'h122 ;
                10'h346 : QQs <= 9'h121 ;
                10'h347 : QQs <= 9'h120 ;
                10'h348 : QQs <= 9'h11F ;
                10'h349 : QQs <= 9'h11E ;
                10'h34A : QQs <= 9'h11D ;
                10'h34B : QQs <= 9'h11C ;
                10'h34C : QQs <= 9'h11A ;
                10'h34D : QQs <= 9'h119 ;
                10'h34E : QQs <= 9'h118 ;
                10'h34F : QQs <= 9'h117 ;
                10'h350 : QQs <= 9'h116 ;
                10'h351 : QQs <= 9'h115 ;
                10'h352 : QQs <= 9'h113 ;
                10'h353 : QQs <= 9'h112 ;
                10'h354 : QQs <= 9'h111 ;
                10'h355 : QQs <= 9'h110 ;
                10'h356 : QQs <= 9'h10F ;
                10'h357 : QQs <= 9'h10E ;
                10'h358 : QQs <= 9'h10C ;
                10'h359 : QQs <= 9'h10B ;
                10'h35A : QQs <= 9'h10A ;
                10'h35B : QQs <= 9'h109 ;
                10'h35C : QQs <= 9'h108 ;
                10'h35D : QQs <= 9'h106 ;
                10'h35E : QQs <= 9'h105 ;
                10'h35F : QQs <= 9'h104 ;
                10'h360 : QQs <= 9'h103 ;
                10'h361 : QQs <= 9'h101 ;
                10'h362 : QQs <= 9'h100 ;
                10'h363 : QQs <= 9'h0FF ;
                10'h364 : QQs <= 9'h0FE ;
                10'h365 : QQs <= 9'h0FC ;
                10'h366 : QQs <= 9'h0FB ;
                10'h367 : QQs <= 9'h0FA ;
                10'h368 : QQs <= 9'h0F9 ;
                10'h369 : QQs <= 9'h0F7 ;
                10'h36A : QQs <= 9'h0F6 ;
                10'h36B : QQs <= 9'h0F5 ;
                10'h36C : QQs <= 9'h0F3 ;
                10'h36D : QQs <= 9'h0F2 ;
                10'h36E : QQs <= 9'h0F1 ;
                10'h36F : QQs <= 9'h0F0 ;
                10'h370 : QQs <= 9'h0EE ;
                10'h371 : QQs <= 9'h0ED ;
                10'h372 : QQs <= 9'h0EC ;
                10'h373 : QQs <= 9'h0EA ;
                10'h374 : QQs <= 9'h0E9 ;
                10'h375 : QQs <= 9'h0E8 ;
                10'h376 : QQs <= 9'h0E6 ;
                10'h377 : QQs <= 9'h0E5 ;
                10'h378 : QQs <= 9'h0E4 ;
                10'h379 : QQs <= 9'h0E2 ;
                10'h37A : QQs <= 9'h0E1 ;
                10'h37B : QQs <= 9'h0E0 ;
                10'h37C : QQs <= 9'h0DE ;
                10'h37D : QQs <= 9'h0DD ;
                10'h37E : QQs <= 9'h0DB ;
                10'h37F : QQs <= 9'h0DA ;
                10'h380 : QQs <= 9'h0D9 ;
                10'h381 : QQs <= 9'h0D7 ;
                10'h382 : QQs <= 9'h0D6 ;
                10'h383 : QQs <= 9'h0D4 ;
                10'h384 : QQs <= 9'h0D3 ;
                10'h385 : QQs <= 9'h0D2 ;
                10'h386 : QQs <= 9'h0D0 ;
                10'h387 : QQs <= 9'h0CF ;
                10'h388 : QQs <= 9'h0CD ;
                10'h389 : QQs <= 9'h0CC ;
                10'h38A : QQs <= 9'h0CB ;
                10'h38B : QQs <= 9'h0C9 ;
                10'h38C : QQs <= 9'h0C8 ;
                10'h38D : QQs <= 9'h0C6 ;
                10'h38E : QQs <= 9'h0C5 ;
                10'h38F : QQs <= 9'h0C3 ;
                10'h390 : QQs <= 9'h0C2 ;
                10'h391 : QQs <= 9'h0C0 ;
                10'h392 : QQs <= 9'h0BF ;
                10'h393 : QQs <= 9'h0BD ;
                10'h394 : QQs <= 9'h0BC ;
                10'h395 : QQs <= 9'h0BA ;
                10'h396 : QQs <= 9'h0B9 ;
                10'h397 : QQs <= 9'h0B7 ;
                10'h398 : QQs <= 9'h0B6 ;
                10'h399 : QQs <= 9'h0B4 ;
                10'h39A : QQs <= 9'h0B3 ;
                10'h39B : QQs <= 9'h0B1 ;
                10'h39C : QQs <= 9'h0B0 ;
                10'h39D : QQs <= 9'h0AE ;
                10'h39E : QQs <= 9'h0AD ;
                10'h39F : QQs <= 9'h0AB ;
                10'h3A0 : QQs <= 9'h0AA ;
                10'h3A1 : QQs <= 9'h0A8 ;
                10'h3A2 : QQs <= 9'h0A7 ;
                10'h3A3 : QQs <= 9'h0A5 ;
                10'h3A4 : QQs <= 9'h0A4 ;
                10'h3A5 : QQs <= 9'h0A2 ;
                10'h3A6 : QQs <= 9'h0A1 ;
                10'h3A7 : QQs <= 9'h09F ;
                10'h3A8 : QQs <= 9'h09D ;
                10'h3A9 : QQs <= 9'h09C ;
                10'h3AA : QQs <= 9'h09A ;
                10'h3AB : QQs <= 9'h099 ;
                10'h3AC : QQs <= 9'h097 ;
                10'h3AD : QQs <= 9'h095 ;
                10'h3AE : QQs <= 9'h094 ;
                10'h3AF : QQs <= 9'h092 ;
                10'h3B0 : QQs <= 9'h091 ;
                10'h3B1 : QQs <= 9'h08F ;
                10'h3B2 : QQs <= 9'h08D ;
                10'h3B3 : QQs <= 9'h08C ;
                10'h3B4 : QQs <= 9'h08A ;
                10'h3B5 : QQs <= 9'h088 ;
                10'h3B6 : QQs <= 9'h087 ;
                10'h3B7 : QQs <= 9'h085 ;
                10'h3B8 : QQs <= 9'h084 ;
                10'h3B9 : QQs <= 9'h082 ;
                10'h3BA : QQs <= 9'h080 ;
                10'h3BB : QQs <= 9'h07F ;
                10'h3BC : QQs <= 9'h07D ;
                10'h3BD : QQs <= 9'h07B ;
                10'h3BE : QQs <= 9'h07A ;
                10'h3BF : QQs <= 9'h078 ;
                10'h3C0 : QQs <= 9'h076 ;
                10'h3C1 : QQs <= 9'h074 ;
                10'h3C2 : QQs <= 9'h073 ;
                10'h3C3 : QQs <= 9'h071 ;
                10'h3C4 : QQs <= 9'h06F ;
                10'h3C5 : QQs <= 9'h06E ;
                10'h3C6 : QQs <= 9'h06C ;
                10'h3C7 : QQs <= 9'h06A ;
                10'h3C8 : QQs <= 9'h068 ;
                10'h3C9 : QQs <= 9'h067 ;
                10'h3CA : QQs <= 9'h065 ;
                10'h3CB : QQs <= 9'h063 ;
                10'h3CC : QQs <= 9'h061 ;
                10'h3CD : QQs <= 9'h060 ;
                10'h3CE : QQs <= 9'h05E ;
                10'h3CF : QQs <= 9'h05C ;
                10'h3D0 : QQs <= 9'h05A ;
                10'h3D1 : QQs <= 9'h059 ;
                10'h3D2 : QQs <= 9'h057 ;
                10'h3D3 : QQs <= 9'h055 ;
                10'h3D4 : QQs <= 9'h053 ;
                10'h3D5 : QQs <= 9'h052 ;
                10'h3D6 : QQs <= 9'h050 ;
                10'h3D7 : QQs <= 9'h04E ;
                10'h3D8 : QQs <= 9'h04C ;
                10'h3D9 : QQs <= 9'h04A ;
                10'h3DA : QQs <= 9'h049 ;
                10'h3DB : QQs <= 9'h047 ;
                10'h3DC : QQs <= 9'h045 ;
                10'h3DD : QQs <= 9'h043 ;
                10'h3DE : QQs <= 9'h041 ;
                10'h3DF : QQs <= 9'h03F ;
                10'h3E0 : QQs <= 9'h03E ;
                10'h3E1 : QQs <= 9'h03C ;
                10'h3E2 : QQs <= 9'h03A ;
                10'h3E3 : QQs <= 9'h038 ;
                10'h3E4 : QQs <= 9'h036 ;
                10'h3E5 : QQs <= 9'h034 ;
                10'h3E6 : QQs <= 9'h032 ;
                10'h3E7 : QQs <= 9'h030 ;
                10'h3E8 : QQs <= 9'h02F ;
                10'h3E9 : QQs <= 9'h02D ;
                10'h3EA : QQs <= 9'h02B ;
                10'h3EB : QQs <= 9'h029 ;
                10'h3EC : QQs <= 9'h027 ;
                10'h3ED : QQs <= 9'h025 ;
                10'h3EE : QQs <= 9'h023 ;
                10'h3EF : QQs <= 9'h021 ;
                10'h3F0 : QQs <= 9'h01F ;
                10'h3F1 : QQs <= 9'h01D ;
                10'h3F2 : QQs <= 9'h01C ;
                10'h3F3 : QQs <= 9'h01A ;
                10'h3F4 : QQs <= 9'h018 ;
                10'h3F5 : QQs <= 9'h016 ;
                10'h3F6 : QQs <= 9'h014 ;
                10'h3F7 : QQs <= 9'h012 ;
                10'h3F8 : QQs <= 9'h010 ;
                10'h3F9 : QQs <= 9'h00E ;
                10'h3FA : QQs <= 9'h00C ;
                10'h3FB : QQs <= 9'h00A ;
                10'h3FC : QQs <= 9'h008 ;
                10'h3FD : QQs <= 9'h006 ;
                10'h3FE : QQs <= 9'h004 ;
                10'h3FF : QQs <= 9'h002 ;
            endcase
        `e
    `r[ 8:0]QQs_D       ;
    `r      CK_EE_DDD   ;
    `ack
        `xar 
        `b
            QQs_D <= 0 ;
            CK_EE_DDD <= 1'b0 ;
        `eelse 
        `b
            CK_EE_DDD <= CK_EE_DD ;
            if( CK_EE_DD ) 
                QQs_D <= QQs ;
        `e
    `a QQs_o = QQs_D ;
    `a B_OUT_DAT_DLYs_o = B_IN_DAT_DLYs_i + C_DAT_DLYs ;
    `a DONE_o = CK_EE_DDD ;
endmodule // SIN_ROM_S11_S11
    `define SIN_ROM_S11_S11
`endif
